library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Entidade que representa a parte operativa do processador MIPS --
entity ParteOperativa is
end entity ParteOperativa;

architecture arch of ParteOperativa is
begin
end arch;
